class xgemac_sequence_item extends uvm_sequence_item;


endclass
