class in_sequence_item extends uvm_sequence_item;


endclass
